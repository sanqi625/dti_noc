`ifndef _PREFIX_
    `define _PREFIX_(x)  Base_``x
`endif