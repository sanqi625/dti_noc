`ifndef _PREFIX_
    `define _PREFIX_(x)  Base_``x
`endif

`ifndef TBU_NUM
    `define TBU_NUM 4
`endif

`ifndef TRANSACTION_MAX_NUM
    `define TRANSACTION_MAX_NUM 8
`endif