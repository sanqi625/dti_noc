package `_PREFIX_(dti_iniu_pack);

    localparam integer unsigned TBU_NUM_WIDTH             = 6;
    localparam integer unsigned AXIS_MAX_DATA_WIDTH       = 160;
    localparam integer unsigned AXIS_DATA_WIDTH           = 80;
    localparam integer unsigned AXIS_KEEP_WIDTH           = AXIS_DATA_WIDTH / 8;
    localparam integer unsigned CUSTOM_DATA_WIDTH         = 80;
    localparam integer unsigned CUSTOM_KEEP_WIDTH         = CUSTOM_DATA_WIDTH / 8;

    typedef enum logic [3:0] {
                              DTI_TBU_CONDIS_REQ = 4'h0,
                              DTI_TBU_TRANS_REQ  = 4'h2
                             } m_msg_type_t;

    typedef enum logic [3:0] {
                              DTI_TBU_CONDIS_ACK   = 4'h0,
                              DTI_TBU_TRANS_FAULT  = 4'h1,
                              DTI_TBU_TRANS_RESP   = 4'h2,
                              DTI_TBU_TRANS_RESPEX = 4'h3
                             } s_msg_type_t;

endpackage