module `_PREFIX_(dti_to_gnpd_conv) 
    import `_PREFIX_(dti_iniu_pack)::*;
    (
    // REQ_data channel
    input   logic                                       req_tvalid                                  ,
    input   logic   [79:0]                              req_tdata                                   ,
    input   logic   [9:0]                               req_tkeep                                   ,
    input   logic                                       req_tlast                                   ,
    input   logic   [5:0]                               req_ttid                                    ,
    output  logic                                       req_tready                                  , //custom rdy
    // RSP_data channel
    output  logic                                       rsp_tvalid                                  ,
    output  logic   [79:0]                              rsp_tdata                                   ,
    output  logic   [9:0]                               rsp_tkeep                                   ,
    output  logic                                       rsp_tlast                                   ,
    output  logic   [5:0]                               rsp_ttid                                    ,
    input   logic                                       rsp_tready                                  , //dti rdy
    // DTI_to_custom
    output logic                                        req_valid                                   ,
    input  logic                                        req_ready                                   ,
    output logic    [89:0]                              req_payload                                 ,
    output logic    [5:0]                               req_srcid                                   ,
    output logic    [5:0]                               req_tgtid                                   ,
    output logic                                        req_qos                                     , //tie1
    output logic                                        req_last                                    ,
    input  logic                                        req_threshold                               , //tie1
    // custom_to_DTI                                                        
    input  logic                                        rsp_valid                                   ,
    output logic                                        rsp_ready                                   ,
    input  logic    [89:0]                              rsp_payload                                 ,
    input  logic    [5:0]                               rsp_srcid                                   ,
    input  logic    [5:0]                               rsp_tgtid                                   ,
    input  logic                                        rsp_qos                                     , //tie 1
    input  logic                                        rsp_last                                    ,
    output logic                                        rsp_threshold                                 //tie 1
    );

    // DTI to custom
    assign req_valid     = req_tvalid;
    assign req_payload   = {req_tdata,req_tkeep};
    assign req_srcid     = req_ttid;
    assign req_tgtid     = 6'd0;
    assign req_qos       = 1'b1; //tie1
    assign req_last      = req_tlast;
    assign req_tready    = req_ready;

    // custom to DTI
    assign rsp_tvalid    = rsp_valid;
    assign rsp_tdata     = rsp_payload[89:10];
    assign rsp_tkeep     = rsp_payload[9:0];
    assign rsp_tlast     = rsp_last;
    assign rsp_ttid      = rsp_srcid;
    assign rsp_threshold = 1'b1; //tie1
    assign rsp_ready     = rsp_tready;

endmodule
