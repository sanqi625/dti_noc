package `_PREFIX_(dti_tniu_pack);

    localparam integer unsigned TBU_NUM_WIDTH             = 6;
    localparam integer unsigned AXIS_DATA_WIDTH           = 80;
    localparam integer unsigned AXIS_KEEP_WIDTH           = AXIS_DATA_WIDTH / 8;
    localparam integer unsigned CUSTOM_DATA_WIDTH         = 80;
    localparam integer unsigned CUSTOM_KEEP_WIDTH         = CUSTOM_DATA_WIDTH / 8;

endpackage